module decoder_4_16(insig, outsig);
	 input [3:0] insig;
	 output [15:0] outsig;
	 reg [15:0] 		outsig;
	 always @ (insig)
		 case(insig)
			 4'b0000: outsig = 16'b0000000000000001;
			 4'b0001: outsig = 16'b0000000000000010;
			 4'b0010: outsig = 16'b0000000000000100;
			 4'b0011: outsig = 16'b0000000000001000;
			 4'b0100: outsig = 16'b0000000000010000;
			 4'b0101: outsig = 16'b0000000000100000;
			 4'b0110: outsig = 16'b0000000001000000;
			 4'b0111: outsig = 16'b0000000010000000;
			 4'b1000: outsig = 16'b0000000100000000;
			 4'b1001: outsig = 16'b0000001000000000;
			 4'b1010: outsig = 16'b0000010000000000;
			 4'b1011: outsig = 16'b0000100000000000;
			 4'b1100: outsig = 16'b0001000000000000;
			 4'b1101: outsig = 16'b0010000000000000;
			 4'b1110: outsig = 16'b0100000000000000;
			 4'b1111: outsig = 16'b1000000000000000;
		 endcase // case (insig)
endmodule // decoder_4_16
